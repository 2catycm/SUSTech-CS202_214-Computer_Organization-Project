module lab1_sw_led_24(
    output[7:0] Minisys_DigitalTubes_NotEnable,
    output[7:0]Minisys_DigitalTube_Shape

    );
    assign Minisys_DigitalTubes_NotEnable = 7'b0000000;
    assign Minisys_DigitalTube_Shape = 7'b0000000;
endmodule

